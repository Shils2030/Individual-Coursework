// Task 3 - 2022
module task3

//Write solution here
		

endmodule
